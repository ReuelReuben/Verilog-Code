module BKA16bit(s,c,a,b,cin);
input [15:0] a,b;
input cin;
output [15:0] s,c;
wire [15:0] p,g;
wire p23,g23,p45,g45,p67,g67,p89,g89,p1011,g1011,p1213,g1213,p1415,g1415;
wire p47,g47,p811,g811,p1215,g1215;
wire p815,g815;

//Pre Processing
Pre b1 (p[0],g[0],a[0],b[0]);
Pre b2 (p[1],g[1],a[1],b[1]);
Pre b3 (p[2],g[2],a[2],b[2]);
Pre b4 (p[3],g[3],a[3],b[3]);
Pre b5 (p[4],g[4],a[4],b[4]);
Pre b6 (p[5],g[5],a[5],b[5]);
Pre b7 (p[6],g[6],a[6],b[6]);
Pre b8 (p[7],g[7],a[7],b[7]);
Pre b9 (p[8],g[8],a[8],b[8]);
Pre b10 (p[9],g[9],a[9],b[9]);
Pre b11 (p[10],g[10],a[10],b[10]);
Pre b12 (p[11],g[11],a[11],b[11]);
Pre b13 (p[12],g[12],a[12],b[12]);
Pre b14 (p[13],g[13],a[13],b[13]);
Pre b15 (p[14],g[14],a[14],b[14]);
Pre b16 (p[15],g[15],a[15],b[15]);

//Stage 1
G b17 (c[0],cin,p[0],g[0]);
G b18 (c[1],c[0],p[1],g[1]);
PG b20 (p23,g23,p[2],g[2],p[3],g[3]);
PG b22 (p45,g45,p[4],g[4],p[5],g[5]);
PG b24 (p67,g67,p[6],g[6],p[7],g[7]);
PG b26 (p89,g89,p[8],g[8],p[9],g[9]);
PG b28 (p1011,g1011,p[10],g[10],p[11],g[11]);
PG b30 (p1213,g1213,p[12],g[12],p[13],g[13]);
PG b32 (p1415,g1415,p[14],g[14],p[15],g[15]);

//Stage 2
G b34 (c[3],c[1],p23,g23);
PG b38 (p47,g47,p45,g45,p67,g67);
PG b42 (p811,g811,p89,g89,p1011,g1011);
PG b46 (p1215,g1215,p1213,g1213,p1415,g1415);

//Stage 3
G b50 (c[7],c[3],p47,g47);
PG b58 (p815,g815,p811,g811,p1215,g1215);

//Stage 4
G b66 (c[15],c[7],p815,g815);

//Stage 5
G b35 (c[2],c[1],p[2],g[2]);
G b67 (c[4],c[3],p[4],g[4]);
G b68 (c[5],c[3],p45,g45);
G b69 (c[6],c[5],p[6],g[6]);
G b70 (c[8],c[7],p[8],g[8]);
G b71 (c[9],c[8],p89,g89);
G b72 (c[10],c[9],p[10],g[10]);
G b73 (c[11],c[7],p811,g811);
G b74 (c[12],c[11],p[12],g[12]);
G b75 (c[13],c[11],p1213,g1213);
G b76 (c[14],c[13],p[14],g[14]);

//Post Processing
xor g1 (s[0],p[0],cin);
xor g2 (s[1],p[1],c[0]);
xor g3 (s[2],p[2],c[1]);
xor g4 (s[3],p[3],c[2]);
xor g5 (s[4],p[4],c[3]);
xor g6 (s[5],p[5],c[4]);
xor g7 (s[6],p[6],c[5]);
xor g8 (s[7],p[7],c[6]);
xor g9 (s[8],p[8],c[7]);
xor g10 (s[9],p[9],c[8]);
xor g11 (s[10],p[10],c[9]);
xor g12 (s[11],p[11],c[10]);
xor g13 (s[12],p[12],c[11]);
xor g14 (s[13],p[13],c[12]);
xor g15 (s[14],p[14],c[13]);
xor g16 (s[15],p[15],c[14]);

endmodule
