module KSA16bit(s,c,a,b,cin);
input [15:0] a,b;
input cin;
output [15:0] s,c;
wire [15:0] p,g;
wire p12,g12,p23,g23,p34,g34,p45,g45,p56,g56,p67,g67,p78,g78,p89,g89,p910,g910,p1011,g1011,p1112,g1112,p1213,g1213,p1314,g1314,p1415,g1415;
wire p14,g14,p25,g25,p36,g36,p47,g47,p58,g58,p69,g69,p710,g710,p811,g811,p912,g912,p1013,g1013,p1114,g1114,p1215,g1215;
wire p18,g18,p29,g29,p310,g310,p411,g411,p512,g512,p613,g613,p714,g714,p815,g815;

//Pre Processing
Pre b1 (p[0],g[0],a[0],b[0]);
Pre b2 (p[1],g[1],a[1],b[1]);
Pre b3 (p[2],g[2],a[2],b[2]);
Pre b4 (p[3],g[3],a[3],b[3]);
Pre b5 (p[4],g[4],a[4],b[4]);
Pre b6 (p[5],g[5],a[5],b[5]);
Pre b7 (p[6],g[6],a[6],b[6]);
Pre b8 (p[7],g[7],a[7],b[7]);
Pre b9 (p[8],g[8],a[8],b[8]);
Pre b10 (p[9],g[9],a[9],b[9]);
Pre b11 (p[10],g[10],a[10],b[10]);
Pre b12 (p[11],g[11],a[11],b[11]);
Pre b13 (p[12],g[12],a[12],b[12]);
Pre b14 (p[13],g[13],a[13],b[13]);
Pre b15 (p[14],g[14],a[14],b[14]);
Pre b16 (p[15],g[15],a[15],b[15]);

//Stage 1
G b17 (c[0],cin,p[0],g[0]);
G b18 (c[1],c[0],p[1],g[1]);
PG b19 (p12,g12,p[1],g[1],p[2],g[2]);
PG b20 (p23,g23,p[2],g[2],p[3],g[3]);
PG b21 (p34,g34,p[3],g[3],p[4],g[4]);
PG b22 (p45,g45,p[4],g[4],p[5],g[5]);
PG b23 (p56,g56,p[5],g[5],p[6],g[6]);
PG b24 (p67,g67,p[6],g[6],p[7],g[7]);
PG b25 (p78,g78,p[7],g[7],p[8],g[8]);
PG b26 (p89,g89,p[8],g[8],p[9],g[9]);
PG b27 (p910,g910,p[9],g[9],p[10],g[10]);
PG b28 (p1011,g1011,p[10],g[10],p[11],g[11]);
PG b29 (p1112,g1112,p[11],g[11],p[12],g[12]);
PG b30 (p1213,g1213,p[12],g[12],p[13],g[13]);
PG b31 (p1314,g1314,p[13],g[13],p[14],g[14]);
PG b32 (p1415,g1415,p[14],g[14],p[15],g[15]);

//Stage 2
G b33 (c[2],c[0],p12,g12);
G b34 (c[3],c[1],p23,g23);
PG b35 (p14,g14,p12,g12,p34,g34);
PG b36 (p25,g25,p23,g23,p45,g45);
PG b37 (p36,g36,p34,g34,p56,g56);
PG b38 (p47,g47,p45,g45,p67,g67);
PG b39 (p58,g58,p56,g56,p78,g78);
PG b40 (p69,g69,p67,g67,p89,g89);
PG b41 (p710,g710,p78,g78,p910,g910);
PG b42 (p811,g811,p89,g89,p1011,g1011);
PG b43 (p912,g912,p910,g910,p1112,g1112);
PG b44 (p1013,g1013,p1011,g1011,p1213,g1213);
PG b45 (p1114,g1114,p1112,g1112,p1314,g1314);
PG b46 (p1215,g1215,p1213,g1213,p1415,g1415);

//Stage 3
G b47 (c[4],c[0],p14,g14);
G b48 (c[5],c[1],p25,g25);
G b49 (c[6],c[2],p36,g36);
G b50 (c[7],c[3],p47,g47);
PG b51 (p18,g18,p14,g14,p58,g58);
PG b52 (p29,g29,p25,g25,p69,g69);
PG b53 (p310,g310,p36,g36,p710,g710);
PG b54 (p411,g411,p47,g47,p811,g811);
PG b55 (p512,g512,p58,g58,p912,g912);
PG b56 (p613,g613,p69,g69,p1013,g1013);
PG b57 (p714,g714,p710,g710,p1114,g1114);
PG b58 (p815,g815,p811,g811,p1215,g1215);

//Stage 4
G b59 (c[8],c[0],p18,g18);
G b60 (c[9],c[1],p29,g29);
G b61 (c[10],c[2],p310,g310);
G b62 (c[11],c[3],p411,g411);
G b63 (c[12],c[4],p512,g512);
G b64 (c[13],c[5],p613,g613);
G b65 (c[14],c[6],p714,g714);
G b66 (c[15],c[7],p815,g815);

//Post Processing
xor g1 (s[0],p[0],cin);
xor g2 (s[1],p[1],c[0]);
xor g3 (s[2],p[2],c[1]);
xor g4 (s[3],p[3],c[2]);
xor g5 (s[4],p[4],c[3]);
xor g6 (s[5],p[5],c[4]);
xor g7 (s[6],p[6],c[5]);
xor g8 (s[7],p[7],c[6]);
xor g9 (s[8],p[8],c[7]);
xor g10 (s[9],p[9],c[8]);
xor g11 (s[10],p[10],c[9]);
xor g12 (s[11],p[11],c[10]);
xor g13 (s[12],p[12],c[11]);
xor g14 (s[13],p[13],c[12]);
xor g15 (s[14],p[14],c[13]);
xor g16 (s[15],p[15],c[14]);

endmodule
